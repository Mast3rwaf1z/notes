library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ex43 is
    port(
        inc : in std_logic;
        dec : in std_logic
    );
end entity ex43;

architecture arch of ex43 is
    signal counter : integer;

begin
    process(inc) is begin
        if rising_edge(inc) then
            counter <= counter + 1;
        end if;
    end process;

    process(dec) is begin
        if counter = 0 then
            counter <= 0;
        elsif rising_edge(dec) then
            counter <= counter - 1;
        end if;
    end process;
end architecture arch;